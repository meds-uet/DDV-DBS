interface add_if;
    logic [3:0] a;
    logic [3:0] b;
    logic [3:0] s;
    logic cin;
    logic cout;
endinterface