interface design_interface(input logic clk_i , reset_i);

logic en_i;
logic [15:0]in1;
logic [15:0]in2;
logic [15:0]sum;


endinterface
