interface add_if;
	logic reset;
	logic clk;
	logic X;
	logic det;
endinterface