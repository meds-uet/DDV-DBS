interface design_interface();

  logic [3:0]in;
  logic [6:0]binary_code;

endinterface
