module design()

endmodule
