// ///////////////Interface Class
interface spi_if;
 
  
  logic clk;
  logic sclk;
  logic newd;
  logic rst;
  logic [11:0] din;
  logic [11:0] dout;
 logic done;
  
  
endinterface