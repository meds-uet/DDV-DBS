module adder_4b(input logic unsigned [3:0] a,b,
                output logic unsigned [4:0] c);


    assign c = a+b;

endmodule
